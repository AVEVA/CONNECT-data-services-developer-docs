[{"type":"Conceptual","source_relative_path":"index.md","output":{".html":{"relative_path":"index.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\qcgc0h23.0wj","hash":"e6SopcHN90OtOA5Dvk1bVw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/SdsStreamExtra.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/SdsStreamExtra.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\p0ckyksw.pe5","hash":"nIJdNG3J3R/64TOSBo9cww=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Reading_Data.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Reading_Data.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\1brxjc0c.1nl","hash":"wb8QUzVgSigHCNPDljHGGA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Quick_Start.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Quick_Start.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\mtvgozid.txz","hash":"Y9CGTiTIDwFnr6eMM5SQnA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataIngress/OMF_Ingress_Specification.md","output":{".html":{"relative_path":"Documentation/DataIngress/OMF_Ingress_Specification.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\oxy0hp0w.3pv","hash":"CHMOs8s9TcoQxUiDvNUAow=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Introducing_SDS.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Introducing_SDS.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\peiasscf.5yc","hash":"cf5siMtagJW0Ik57pR6CqQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_ClientRole.md","output":{".html":{"relative_path":"Documentation/Management/Account_ClientRole.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\zxzdyrwy.y4q","hash":"t6q6WZhQVlTIofOy04UJxA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_Namespace.md","output":{".html":{"relative_path":"Documentation/Management/Account_Namespace.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\2rnhbot2.53e","hash":"UTlP2Vykxtd5qpJrLzrg+g=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_NamespaceTier.md","output":{".html":{"relative_path":"Documentation/Management/Account_NamespaceTier.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\cltvytv0.kaz","hash":"2gtPuSZNa3RbT2F7h6cq0Q=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_Role.md","output":{".html":{"relative_path":"Documentation/Management/Account_Role.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\wucf3g4r.3dj","hash":"juzdPf1x7FvQVac8TfPwQA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_RootAccessControl.md","output":{".html":{"relative_path":"Documentation/Management/Account_RootAccessControl.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\3qx3mol5.4zu","hash":"w/pYza1vtqk99SHJ9jDSSg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_ServiceBlog.md","output":{".html":{"relative_path":"Documentation/Management/Account_ServiceBlog.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\q3ypigvq.skc","hash":"Qn+emR3cTkPVxoGkOtGW6g=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_Tenant.md","output":{".html":{"relative_path":"Documentation/Management/Account_Tenant.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\c0ojhbao.xz4","hash":"+877gbuh5r7JNGjZiWKqCQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_TenantFeatureState.md","output":{".html":{"relative_path":"Documentation/Management/Account_TenantFeatureState.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\sdixgmqs.xo5","hash":"a+VvYEfWYVwNEOVT7OQVyA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Account_UserRole.md","output":{".html":{"relative_path":"Documentation/Management/Account_UserRole.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\454uythr.n0y","hash":"9cnox9UNrlC2qy1xb8PEew=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/SDS_Types.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/SDS_Types.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ryrdhm2v.fmx","hash":"bONXtbqnSGv//OnWXa9PLQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/SDS_Streams.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/SDS_Streams.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\adpqlekh.33b","hash":"p3qWwspNSM0yPNfgdAQgTg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Filter_Expressions_Metadata.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Filter_Expressions_Metadata.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\s25oi1o0.qsj","hash":"VY180p/67hHFYi9bFDXZKA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Management/Management_Overview.md","output":{".html":{"relative_path":"Documentation/Management/Management_Overview.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\evxee1kx.xww","hash":"pnV3jJM4cn0sW5rBk4+KEg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Units_of_Measure.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Units_of_Measure.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\zhcfpuez.rr5","hash":"TeuVJ6+cy+pK5odRSjE4cw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Searching.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Searching.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\yeedbkng.gt4","hash":"djlp6s2C+5JcXQrwmHPFQQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_HybridClient.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_HybridClient.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\lidya4um.1r2","hash":"LZVGmlM5ODfzQzWEtyIfsQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_Client.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_Client.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ova4g1xo.5dj","hash":"Mbobt+tuzp7E1C0nJySAUg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_ClientCredentialClient.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_ClientCredentialClient.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\11viehim.doi","hash":"5akqakeYkPMpnLBAYOMpHA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_IdentityProvider.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_IdentityProvider.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ans3odwz.b2d","hash":"f6wQEl0gm1IBQLEAekFLFw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_ImplicitClient.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_ImplicitClient.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\1bem1osf.pmo","hash":"cdHGW6Df1zDSbiHLnGAJdw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_Invitation.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_Invitation.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\w50ysdgp.ogl","hash":"qIMCH19bCbbk917UiRYKjA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_Secret.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_Secret.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\d1fjaqhd.n0y","hash":"kq2aEn2uNFuP+uCKCWzfrw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_User.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_User.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\041stolz.rf4","hash":"kd4zZ1B3evp9HeC8XPfwsQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/table_format.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/table_format.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\uwj14y1r.oe5","hash":"efvLG8Vhs8OwUNbpgRPZBw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Writing_Data.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Writing_Data.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\mlcbmgmt.eyt","hash":"Iy94rithUQ+S6Cl4NOv1nw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Writing_Data_API.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Writing_Data_API.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ol2qt0mb.q5u","hash":"9O+VAfcRiBS55cisL9BBEA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/support.md","output":{".html":{"relative_path":"Documentation/support.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\qb40wese.wi0","hash":"t240QA7r9BQkIfAFuozcUg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Access_Control.md","output":{".html":{"relative_path":"Documentation/Access_Control.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\jcmmur3w.wae","hash":"AmVlLenh1LK8lAiEhHFrOQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/OSIsoft_Cloud_Services.md","output":{".html":{"relative_path":"Documentation/OSIsoft_Cloud_Services.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\nktdwvqn.314","hash":"EVhppEk6k02bYucEleHm7Q=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataViews/DataViews_Overview.md","output":{".html":{"relative_path":"Documentation/DataViews/DataViews_Overview.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\xtvcr55z.lhl","hash":"GU2dqGNr5CjlvbqzVu0tdw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataViews/DataViews_API.md","output":{".html":{"relative_path":"Documentation/DataViews/DataViews_API.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\klij3wkv.swk","hash":"ibYGUc2YGl0A6/CZ2qRPQw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Data_Store_and_SDS.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Data_Store_and_SDS.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\0ol5kgd3.lld","hash":"XRh/RFnFW0rcQlIcQ0xCwg=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Identity_Overview.md","output":{".html":{"relative_path":"Documentation/Identity/Identity_Overview.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\i1zp130h.ru3","hash":"TFCOl2zjUmUXo3OUqy2uZw=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/Identity/Consent.md","output":{".html":{"relative_path":"Documentation/Identity/Consent.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\h4etf5ob.id4","hash":"cvIc3AiaHXR48E2Z4P6hcQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataIngress/OMF_Ingress_Subscriptions.md","output":{".html":{"relative_path":"Documentation/DataIngress/OMF_Ingress_Subscriptions.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\riyn3jgc.bdo","hash":"IbVcyji4rdFl3HUuURLqoA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Filter_Expressions.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Filter_Expressions.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\31zrs14w.qbj","hash":"fLVEqWJMTJ6kmjANBSGUaA=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/indexes.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/indexes.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ji3yjedc.2c2","hash":"FKaB5cSqlsvSl58bCcDiLQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataIngress/OMF_Ingress_to_OCS.md","output":{".html":{"relative_path":"Documentation/DataIngress/OMF_Ingress_to_OCS.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\sialpbml.zvi","hash":"Xv+2HESE87BZA6HWKCsuhQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataIngress/OMF_Ingress_Topics.md","output":{".html":{"relative_path":"Documentation/DataIngress/OMF_Ingress_Topics.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\fzcbmjo2.5r4","hash":"B6EMjzqP7qbWACSqHN/1lQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/DataIngress/Data_Ingress.md","output":{".html":{"relative_path":"Documentation/DataIngress/Data_Ingress.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\upcx4f3p.4o4","hash":"Ks+EYXCArkWV8CWl+t65JQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/samples.md","output":{".html":{"relative_path":"Documentation/samples.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\pi0uch1c.0nx","hash":"iofRCtN5xnz3bXpKiWc2FQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Reading_Data_API.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Reading_Data_API.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\ms10zvzn.un4","hash":"gpOnCqdBeExjvAlZin3XNQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/SDS_Views.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/SDS_Views.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\hp4focde.gum","hash":"CTfxN7ugjh9Fy0qpF7QBQQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"Documentation/SequentialDataStore/Compression.md","output":{".html":{"relative_path":"Documentation/SequentialDataStore/Compression.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\qzwsh0pf.lpw","hash":"3ED2cyC1dvFA/B8uz60JVg=="}},"is_incremental":true,"version":""},{"type":"Toc","source_relative_path":"Documentation/toc.yml","output":{".html":{"relative_path":"Documentation/toc.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\vgmgefgc.2tm","hash":"CTj5FQpcrNdvnPaezZAhkA=="}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/Add_Button.png","output":{"resource":{"relative_path":"Documentation/images/Add_Button.png","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/Add_Button.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/Acquire_Token.png","output":{"resource":{"relative_path":"Documentation/images/Acquire_Token.png","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/Acquire_Token.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous1.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous1.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous1.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsSimpleDiscrete.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsSimpleDiscrete.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsSimpleDiscrete.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsComplexType.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsComplexType.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsComplexType.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/atlas_icon.png","output":{"resource":{"relative_path":"Documentation/images/atlas_icon.png","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/atlas_icon.png"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/Acquire_Client_Key.png","output":{"resource":{"relative_path":"Documentation/images/Acquire_Client_Key.png","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/Acquire_Client_Key.png"}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"toc.yml","output":{".html":{"relative_path":"toc.html","link_to_path":"C:\\agent\\_work\\5\\s\\obj\\.cache\\build\\libos1zg.nfx\\qboj0nlr.y2x","hash":"crXFTLtj6FStiF2rM/zh1g=="}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsSimpleType.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsSimpleType.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsSimpleType.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous2.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous2.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsSimpleStepwiseContinuous2.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsSimpleContinuous.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsSimpleContinuous.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsSimpleContinuous.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/QiDataBehaviorsComplexTypeWithBehavior.PNG","output":{"resource":{"relative_path":"Documentation/images/QiDataBehaviorsComplexTypeWithBehavior.PNG","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/QiDataBehaviorsComplexTypeWithBehavior.PNG"}},"is_incremental":false,"version":""},{"type":"Resource","source_relative_path":"Documentation/images/Containers_1A.png","output":{"resource":{"relative_path":"Documentation/images/Containers_1A.png","link_to_path":"C:\\agent\\_work\\5\\s/Documentation/images/Containers_1A.png"}},"is_incremental":false,"version":""}]